
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity SHR is
  Port ( 
    X: in unsigned(31 downto 0);
    Result : out unsigned(31 downto 0)
    );
end SHR;

architecture SHR of SHR is

begin


end SHR;
